-- qsys0.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity qsys0 is
	port (
		clk_clk       : in    std_logic                     := '0';             --   clk.clk
		gpio_export   : inout std_logic_vector(31 downto 0) := (others => '0'); --  gpio.export
		jtag_tms      : in    std_logic                     := '0';             --  jtag.tms
		jtag_tdi      : in    std_logic                     := '0';             --      .tdi
		jtag_tdo      : out   std_logic;                                        --      .tdo
		jtag_tck      : in    std_logic                     := '0';             --      .tck
		reset_reset_n : in    std_logic                     := '0';             -- reset.reset_n
		uart_rxd      : in    std_logic                     := '0';             --  uart.rxd
		uart_txd      : out   std_logic                                         --      .txd
	);
end entity qsys0;

architecture rtl of qsys0 is
	component VexRiscvAvalon is
		generic (
			C_RESET_VECTOR     : std_logic_vector(31 downto 0) := "00000000000000000000000000010000";
			C_EXCEPTION_VECTOR : std_logic_vector(31 downto 0) := "00000000000000000000000000100000";
			C_IO_BEGIN         : std_logic_vector(31 downto 0) := "10000000000000000000000000000000";
			C_IO_END           : std_logic_vector(31 downto 0) := "11111111111111111111111111111111";
			CORE_CONFIG        : natural                       := 1
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			jtag_tms                 : in  std_logic                     := 'X';             -- export
			jtag_tdi                 : in  std_logic                     := 'X';             -- export
			jtag_tdo                 : out std_logic;                                        -- export
			jtag_tck                 : in  std_logic                     := 'X';             -- export
			iBusAvalon_address       : out std_logic_vector(31 downto 0);                    -- address
			iBusAvalon_read          : out std_logic;                                        -- read
			iBusAvalon_waitRequestn  : in  std_logic                     := 'X';             -- waitrequest_n
			iBusAvalon_response      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			iBusAvalon_readDataValid : in  std_logic                     := 'X';             -- readdatavalid
			iBusAvalon_readData      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dBusAvalon_address       : out std_logic_vector(31 downto 0);                    -- address
			dBusAvalon_read          : out std_logic;                                        -- read
			dBusAvalon_write         : out std_logic;                                        -- write
			dBusAvalon_waitRequestn  : in  std_logic                     := 'X';             -- waitrequest_n
			dBusAvalon_byteEnable    : out std_logic_vector(3 downto 0);                     -- byteenable
			dBusAvalon_writeData     : out std_logic_vector(31 downto 0);                    -- writedata
			dBusAvalon_response      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			dBusAvalon_readDataValid : in  std_logic                     := 'X';             -- readdatavalid
			dBusAvalon_readData      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ic_avalon_address        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			ic_avalon_write          : in  std_logic                     := 'X';             -- write
			ic_avalon_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ic_avalon_read           : in  std_logic                     := 'X';             -- read
			ic_avalon_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			ic_avalon_readdatavalid  : out std_logic;                                        -- readdatavalid
			ic_avalon_waitrequest    : out std_logic;                                        -- waitrequest
			irq_source               : in  std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component VexRiscvAvalon;

	component qsys0_onchip_memory2_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component qsys0_onchip_memory2_0;

	component qsys0_pio_0 is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component qsys0_pio_0;

	component qsys0_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component qsys0_uart_0;

	component qsys0_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			VexRiscvAvalon_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			VexRiscvAvalon_0_data_bus_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			VexRiscvAvalon_0_data_bus_waitrequest              : out std_logic;                                        -- waitrequest
			VexRiscvAvalon_0_data_bus_byteenable               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			VexRiscvAvalon_0_data_bus_read                     : in  std_logic                     := 'X';             -- read
			VexRiscvAvalon_0_data_bus_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			VexRiscvAvalon_0_data_bus_readdatavalid            : out std_logic;                                        -- readdatavalid
			VexRiscvAvalon_0_data_bus_write                    : in  std_logic                     := 'X';             -- write
			VexRiscvAvalon_0_data_bus_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			VexRiscvAvalon_0_data_bus_response                 : out std_logic_vector(1 downto 0);                     -- response
			onchip_memory2_0_s2_address                        : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s2_write                          : out std_logic;                                        -- write
			onchip_memory2_0_s2_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s2_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s2_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s2_chipselect                     : out std_logic;                                        -- chipselect
			onchip_memory2_0_s2_clken                          : out std_logic;                                        -- clken
			pio_0_s1_address                                   : out std_logic_vector(2 downto 0);                     -- address
			pio_0_s1_write                                     : out std_logic;                                        -- write
			pio_0_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_0_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_s1_chipselect                                : out std_logic;                                        -- chipselect
			uart_0_s1_address                                  : out std_logic_vector(2 downto 0);                     -- address
			uart_0_s1_write                                    : out std_logic;                                        -- write
			uart_0_s1_read                                     : out std_logic;                                        -- read
			uart_0_s1_readdata                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_0_s1_writedata                                : out std_logic_vector(15 downto 0);                    -- writedata
			uart_0_s1_begintransfer                            : out std_logic;                                        -- begintransfer
			uart_0_s1_chipselect                               : out std_logic;                                        -- chipselect
			VexRiscvAvalon_0_irq_controller_address            : out std_logic_vector(3 downto 0);                     -- address
			VexRiscvAvalon_0_irq_controller_write              : out std_logic;                                        -- write
			VexRiscvAvalon_0_irq_controller_read               : out std_logic;                                        -- read
			VexRiscvAvalon_0_irq_controller_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			VexRiscvAvalon_0_irq_controller_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			VexRiscvAvalon_0_irq_controller_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			VexRiscvAvalon_0_irq_controller_waitrequest        : in  std_logic                     := 'X'              -- waitrequest
		);
	end component qsys0_mm_interconnect_0;

	component qsys0_mm_interconnect_1 is
		port (
			clk_0_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			VexRiscvAvalon_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			VexRiscvAvalon_0_instruction_bus_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			VexRiscvAvalon_0_instruction_bus_waitrequest       : out std_logic;                                        -- waitrequest
			VexRiscvAvalon_0_instruction_bus_read              : in  std_logic                     := 'X';             -- read
			VexRiscvAvalon_0_instruction_bus_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			VexRiscvAvalon_0_instruction_bus_readdatavalid     : out std_logic;                                        -- readdatavalid
			VexRiscvAvalon_0_instruction_bus_response          : out std_logic_vector(1 downto 0);                     -- response
			onchip_memory2_0_s1_address                        : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s1_write                          : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                     : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                     : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                          : out std_logic                                         -- clken
		);
	end component qsys0_mm_interconnect_1;

	component qsys0_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component qsys0_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal mm_interconnect_0_vexriscvavalon_0_data_bus_waitrequest         : std_logic;                     -- mm_interconnect_0:VexRiscvAvalon_0_data_bus_waitrequest -> mm_interconnect_0_vexriscvavalon_0_data_bus_waitrequest:in
	signal vexriscvavalon_0_data_bus_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:VexRiscvAvalon_0_data_bus_readdata -> VexRiscvAvalon_0:dBusAvalon_readData
	signal vexriscvavalon_0_data_bus_address                               : std_logic_vector(31 downto 0); -- VexRiscvAvalon_0:dBusAvalon_address -> mm_interconnect_0:VexRiscvAvalon_0_data_bus_address
	signal vexriscvavalon_0_data_bus_read                                  : std_logic;                     -- VexRiscvAvalon_0:dBusAvalon_read -> mm_interconnect_0:VexRiscvAvalon_0_data_bus_read
	signal vexriscvavalon_0_data_bus_byteenable                            : std_logic_vector(3 downto 0);  -- VexRiscvAvalon_0:dBusAvalon_byteEnable -> mm_interconnect_0:VexRiscvAvalon_0_data_bus_byteenable
	signal vexriscvavalon_0_data_bus_readdatavalid                         : std_logic;                     -- mm_interconnect_0:VexRiscvAvalon_0_data_bus_readdatavalid -> VexRiscvAvalon_0:dBusAvalon_readDataValid
	signal vexriscvavalon_0_data_bus_response                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:VexRiscvAvalon_0_data_bus_response -> VexRiscvAvalon_0:dBusAvalon_response
	signal vexriscvavalon_0_data_bus_write                                 : std_logic;                     -- VexRiscvAvalon_0:dBusAvalon_write -> mm_interconnect_0:VexRiscvAvalon_0_data_bus_write
	signal vexriscvavalon_0_data_bus_writedata                             : std_logic_vector(31 downto 0); -- VexRiscvAvalon_0:dBusAvalon_writeData -> mm_interconnect_0:VexRiscvAvalon_0_data_bus_writedata
	signal mm_interconnect_0_vexriscvavalon_0_irq_controller_readdata      : std_logic_vector(31 downto 0); -- VexRiscvAvalon_0:ic_avalon_readdata -> mm_interconnect_0:VexRiscvAvalon_0_irq_controller_readdata
	signal mm_interconnect_0_vexriscvavalon_0_irq_controller_waitrequest   : std_logic;                     -- VexRiscvAvalon_0:ic_avalon_waitrequest -> mm_interconnect_0:VexRiscvAvalon_0_irq_controller_waitrequest
	signal mm_interconnect_0_vexriscvavalon_0_irq_controller_address       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:VexRiscvAvalon_0_irq_controller_address -> VexRiscvAvalon_0:ic_avalon_address
	signal mm_interconnect_0_vexriscvavalon_0_irq_controller_read          : std_logic;                     -- mm_interconnect_0:VexRiscvAvalon_0_irq_controller_read -> VexRiscvAvalon_0:ic_avalon_read
	signal mm_interconnect_0_vexriscvavalon_0_irq_controller_readdatavalid : std_logic;                     -- VexRiscvAvalon_0:ic_avalon_readdatavalid -> mm_interconnect_0:VexRiscvAvalon_0_irq_controller_readdatavalid
	signal mm_interconnect_0_vexriscvavalon_0_irq_controller_write         : std_logic;                     -- mm_interconnect_0:VexRiscvAvalon_0_irq_controller_write -> VexRiscvAvalon_0:ic_avalon_write
	signal mm_interconnect_0_vexriscvavalon_0_irq_controller_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:VexRiscvAvalon_0_irq_controller_writedata -> VexRiscvAvalon_0:ic_avalon_writedata
	signal mm_interconnect_0_pio_0_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	signal mm_interconnect_0_pio_0_s1_readdata                             : std_logic_vector(31 downto 0); -- pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	signal mm_interconnect_0_pio_0_s1_address                              : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pio_0_s1_address -> pio_0:address
	signal mm_interconnect_0_pio_0_s1_write                                : std_logic;                     -- mm_interconnect_0:pio_0_s1_write -> mm_interconnect_0_pio_0_s1_write:in
	signal mm_interconnect_0_pio_0_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	signal mm_interconnect_0_uart_0_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	signal mm_interconnect_0_uart_0_s1_readdata                            : std_logic_vector(15 downto 0); -- uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	signal mm_interconnect_0_uart_0_s1_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_0_s1_address -> uart_0:address
	signal mm_interconnect_0_uart_0_s1_read                                : std_logic;                     -- mm_interconnect_0:uart_0_s1_read -> mm_interconnect_0_uart_0_s1_read:in
	signal mm_interconnect_0_uart_0_s1_begintransfer                       : std_logic;                     -- mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	signal mm_interconnect_0_uart_0_s1_write                               : std_logic;                     -- mm_interconnect_0:uart_0_s1_write -> mm_interconnect_0_uart_0_s1_write:in
	signal mm_interconnect_0_uart_0_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s2_chipselect                : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	signal mm_interconnect_0_onchip_memory2_0_s2_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	signal mm_interconnect_0_onchip_memory2_0_s2_address                   : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	signal mm_interconnect_0_onchip_memory2_0_s2_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	signal mm_interconnect_0_onchip_memory2_0_s2_write                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	signal mm_interconnect_0_onchip_memory2_0_s2_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	signal mm_interconnect_0_onchip_memory2_0_s2_clken                     : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	signal mm_interconnect_1_vexriscvavalon_0_instruction_bus_waitrequest  : std_logic;                     -- mm_interconnect_1:VexRiscvAvalon_0_instruction_bus_waitrequest -> mm_interconnect_1_vexriscvavalon_0_instruction_bus_waitrequest:in
	signal vexriscvavalon_0_instruction_bus_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_1:VexRiscvAvalon_0_instruction_bus_readdata -> VexRiscvAvalon_0:iBusAvalon_readData
	signal vexriscvavalon_0_instruction_bus_address                        : std_logic_vector(31 downto 0); -- VexRiscvAvalon_0:iBusAvalon_address -> mm_interconnect_1:VexRiscvAvalon_0_instruction_bus_address
	signal vexriscvavalon_0_instruction_bus_read                           : std_logic;                     -- VexRiscvAvalon_0:iBusAvalon_read -> mm_interconnect_1:VexRiscvAvalon_0_instruction_bus_read
	signal vexriscvavalon_0_instruction_bus_readdatavalid                  : std_logic;                     -- mm_interconnect_1:VexRiscvAvalon_0_instruction_bus_readdatavalid -> VexRiscvAvalon_0:iBusAvalon_readDataValid
	signal vexriscvavalon_0_instruction_bus_response                       : std_logic_vector(1 downto 0);  -- mm_interconnect_1:VexRiscvAvalon_0_instruction_bus_response -> VexRiscvAvalon_0:iBusAvalon_response
	signal mm_interconnect_1_onchip_memory2_0_s1_chipselect                : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_1_onchip_memory2_0_s1_readdata                  : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	signal mm_interconnect_1_onchip_memory2_0_s1_address                   : std_logic_vector(12 downto 0); -- mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_1_onchip_memory2_0_s1_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_1_onchip_memory2_0_s1_write                     : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_1_onchip_memory2_0_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_1_onchip_memory2_0_s1_clken                     : std_logic;                     -- mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- uart_0:irq -> irq_mapper:receiver0_irq
	signal vexriscvavalon_0_interrupt_receiver_irq                         : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> VexRiscvAvalon_0:irq_source
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [VexRiscvAvalon_0:reset, irq_mapper:reset, mm_interconnect_0:VexRiscvAvalon_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:VexRiscvAvalon_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, onchip_memory2_0:reset2, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_0:reset_req2, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal vexriscvavalon_0_data_bus_inv                                   : std_logic;                     -- mm_interconnect_0_vexriscvavalon_0_data_bus_waitrequest:inv -> VexRiscvAvalon_0:dBusAvalon_waitRequestn
	signal mm_interconnect_0_pio_0_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_pio_0_s1_write:inv -> pio_0:write_n
	signal mm_interconnect_0_uart_0_s1_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_uart_0_s1_read:inv -> uart_0:read_n
	signal mm_interconnect_0_uart_0_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_uart_0_s1_write:inv -> uart_0:write_n
	signal vexriscvavalon_0_instruction_bus_inv                            : std_logic;                     -- mm_interconnect_1_vexriscvavalon_0_instruction_bus_waitrequest:inv -> VexRiscvAvalon_0:iBusAvalon_waitRequestn
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [pio_0:reset_n, uart_0:reset_n]

begin

	vexriscvavalon_0 : component VexRiscvAvalon
		generic map (
			C_RESET_VECTOR     => "00000000000000000000000000010000",
			C_EXCEPTION_VECTOR => "00000000000000000000000000100000",
			C_IO_BEGIN         => "00000000000000010000000000000000",
			C_IO_END           => "00000000000000011111111111111111",
			CORE_CONFIG        => 1
		)
		port map (
			clk                      => clk_clk,                                                         --              clock.clk
			reset                    => rst_controller_reset_out_reset,                                  --              reset.reset
			jtag_tms                 => jtag_tms,                                                        --               jtag.export
			jtag_tdi                 => jtag_tdi,                                                        --                   .export
			jtag_tdo                 => jtag_tdo,                                                        --                   .export
			jtag_tck                 => jtag_tck,                                                        --                   .export
			iBusAvalon_address       => vexriscvavalon_0_instruction_bus_address,                        --    instruction_bus.address
			iBusAvalon_read          => vexriscvavalon_0_instruction_bus_read,                           --                   .read
			iBusAvalon_waitRequestn  => vexriscvavalon_0_instruction_bus_inv,                            --                   .waitrequest_n
			iBusAvalon_response      => vexriscvavalon_0_instruction_bus_response,                       --                   .response
			iBusAvalon_readDataValid => vexriscvavalon_0_instruction_bus_readdatavalid,                  --                   .readdatavalid
			iBusAvalon_readData      => vexriscvavalon_0_instruction_bus_readdata,                       --                   .readdata
			dBusAvalon_address       => vexriscvavalon_0_data_bus_address,                               --           data_bus.address
			dBusAvalon_read          => vexriscvavalon_0_data_bus_read,                                  --                   .read
			dBusAvalon_write         => vexriscvavalon_0_data_bus_write,                                 --                   .write
			dBusAvalon_waitRequestn  => vexriscvavalon_0_data_bus_inv,                                   --                   .waitrequest_n
			dBusAvalon_byteEnable    => vexriscvavalon_0_data_bus_byteenable,                            --                   .byteenable
			dBusAvalon_writeData     => vexriscvavalon_0_data_bus_writedata,                             --                   .writedata
			dBusAvalon_response      => vexriscvavalon_0_data_bus_response,                              --                   .response
			dBusAvalon_readDataValid => vexriscvavalon_0_data_bus_readdatavalid,                         --                   .readdatavalid
			dBusAvalon_readData      => vexriscvavalon_0_data_bus_readdata,                              --                   .readdata
			ic_avalon_address        => mm_interconnect_0_vexriscvavalon_0_irq_controller_address,       --     irq_controller.address
			ic_avalon_write          => mm_interconnect_0_vexriscvavalon_0_irq_controller_write,         --                   .write
			ic_avalon_writedata      => mm_interconnect_0_vexriscvavalon_0_irq_controller_writedata,     --                   .writedata
			ic_avalon_read           => mm_interconnect_0_vexriscvavalon_0_irq_controller_read,          --                   .read
			ic_avalon_readdata       => mm_interconnect_0_vexriscvavalon_0_irq_controller_readdata,      --                   .readdata
			ic_avalon_readdatavalid  => mm_interconnect_0_vexriscvavalon_0_irq_controller_readdatavalid, --                   .readdatavalid
			ic_avalon_waitrequest    => mm_interconnect_0_vexriscvavalon_0_irq_controller_waitrequest,   --                   .waitrequest
			irq_source               => vexriscvavalon_0_interrupt_receiver_irq                          -- interrupt_receiver.irq
		);

	onchip_memory2_0 : component qsys0_onchip_memory2_0
		port map (
			clk         => clk_clk,                                          --   clk1.clk
			address     => mm_interconnect_1_onchip_memory2_0_s1_address,    --     s1.address
			clken       => mm_interconnect_1_onchip_memory2_0_s1_clken,      --       .clken
			chipselect  => mm_interconnect_1_onchip_memory2_0_s1_chipselect, --       .chipselect
			write       => mm_interconnect_1_onchip_memory2_0_s1_write,      --       .write
			readdata    => mm_interconnect_1_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_1_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_1_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,               --       .reset_req
			address2    => mm_interconnect_0_onchip_memory2_0_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_onchip_memory2_0_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_onchip_memory2_0_s2_clken,      --       .clken
			write2      => mm_interconnect_0_onchip_memory2_0_s2_write,      --       .write
			readdata2   => mm_interconnect_0_onchip_memory2_0_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_onchip_memory2_0_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_onchip_memory2_0_s2_byteenable, --       .byteenable
			clk2        => clk_clk,                                          --   clk2.clk
			reset2      => rst_controller_reset_out_reset,                   -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze      => '0'                                               -- (terminated)
		);

	pio_0 : component qsys0_pio_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_0_s1_readdata,        --                    .readdata
			bidir_port => gpio_export                                 -- external_connection.export
		);

	uart_0 : component qsys0_uart_0
		port map (
			clk           => clk_clk,                                     --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address       => mm_interconnect_0_uart_0_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_0_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_0_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_0_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_0_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_0_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_0_s1_readdata,        --                    .readdata
			rxd           => uart_rxd,                                    -- external_connection.export
			txd           => uart_txd,                                    --                    .export
			irq           => irq_mapper_receiver0_irq                     --                 irq.irq
		);

	mm_interconnect_0 : component qsys0_mm_interconnect_0
		port map (
			clk_0_clk_clk                                      => clk_clk,                                                         --                                    clk_0_clk.clk
			VexRiscvAvalon_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                  -- VexRiscvAvalon_0_reset_reset_bridge_in_reset.reset
			VexRiscvAvalon_0_data_bus_address                  => vexriscvavalon_0_data_bus_address,                               --                    VexRiscvAvalon_0_data_bus.address
			VexRiscvAvalon_0_data_bus_waitrequest              => mm_interconnect_0_vexriscvavalon_0_data_bus_waitrequest,         --                                             .waitrequest
			VexRiscvAvalon_0_data_bus_byteenable               => vexriscvavalon_0_data_bus_byteenable,                            --                                             .byteenable
			VexRiscvAvalon_0_data_bus_read                     => vexriscvavalon_0_data_bus_read,                                  --                                             .read
			VexRiscvAvalon_0_data_bus_readdata                 => vexriscvavalon_0_data_bus_readdata,                              --                                             .readdata
			VexRiscvAvalon_0_data_bus_readdatavalid            => vexriscvavalon_0_data_bus_readdatavalid,                         --                                             .readdatavalid
			VexRiscvAvalon_0_data_bus_write                    => vexriscvavalon_0_data_bus_write,                                 --                                             .write
			VexRiscvAvalon_0_data_bus_writedata                => vexriscvavalon_0_data_bus_writedata,                             --                                             .writedata
			VexRiscvAvalon_0_data_bus_response                 => vexriscvavalon_0_data_bus_response,                              --                                             .response
			onchip_memory2_0_s2_address                        => mm_interconnect_0_onchip_memory2_0_s2_address,                   --                          onchip_memory2_0_s2.address
			onchip_memory2_0_s2_write                          => mm_interconnect_0_onchip_memory2_0_s2_write,                     --                                             .write
			onchip_memory2_0_s2_readdata                       => mm_interconnect_0_onchip_memory2_0_s2_readdata,                  --                                             .readdata
			onchip_memory2_0_s2_writedata                      => mm_interconnect_0_onchip_memory2_0_s2_writedata,                 --                                             .writedata
			onchip_memory2_0_s2_byteenable                     => mm_interconnect_0_onchip_memory2_0_s2_byteenable,                --                                             .byteenable
			onchip_memory2_0_s2_chipselect                     => mm_interconnect_0_onchip_memory2_0_s2_chipselect,                --                                             .chipselect
			onchip_memory2_0_s2_clken                          => mm_interconnect_0_onchip_memory2_0_s2_clken,                     --                                             .clken
			pio_0_s1_address                                   => mm_interconnect_0_pio_0_s1_address,                              --                                     pio_0_s1.address
			pio_0_s1_write                                     => mm_interconnect_0_pio_0_s1_write,                                --                                             .write
			pio_0_s1_readdata                                  => mm_interconnect_0_pio_0_s1_readdata,                             --                                             .readdata
			pio_0_s1_writedata                                 => mm_interconnect_0_pio_0_s1_writedata,                            --                                             .writedata
			pio_0_s1_chipselect                                => mm_interconnect_0_pio_0_s1_chipselect,                           --                                             .chipselect
			uart_0_s1_address                                  => mm_interconnect_0_uart_0_s1_address,                             --                                    uart_0_s1.address
			uart_0_s1_write                                    => mm_interconnect_0_uart_0_s1_write,                               --                                             .write
			uart_0_s1_read                                     => mm_interconnect_0_uart_0_s1_read,                                --                                             .read
			uart_0_s1_readdata                                 => mm_interconnect_0_uart_0_s1_readdata,                            --                                             .readdata
			uart_0_s1_writedata                                => mm_interconnect_0_uart_0_s1_writedata,                           --                                             .writedata
			uart_0_s1_begintransfer                            => mm_interconnect_0_uart_0_s1_begintransfer,                       --                                             .begintransfer
			uart_0_s1_chipselect                               => mm_interconnect_0_uart_0_s1_chipselect,                          --                                             .chipselect
			VexRiscvAvalon_0_irq_controller_address            => mm_interconnect_0_vexriscvavalon_0_irq_controller_address,       --              VexRiscvAvalon_0_irq_controller.address
			VexRiscvAvalon_0_irq_controller_write              => mm_interconnect_0_vexriscvavalon_0_irq_controller_write,         --                                             .write
			VexRiscvAvalon_0_irq_controller_read               => mm_interconnect_0_vexriscvavalon_0_irq_controller_read,          --                                             .read
			VexRiscvAvalon_0_irq_controller_readdata           => mm_interconnect_0_vexriscvavalon_0_irq_controller_readdata,      --                                             .readdata
			VexRiscvAvalon_0_irq_controller_writedata          => mm_interconnect_0_vexriscvavalon_0_irq_controller_writedata,     --                                             .writedata
			VexRiscvAvalon_0_irq_controller_readdatavalid      => mm_interconnect_0_vexriscvavalon_0_irq_controller_readdatavalid, --                                             .readdatavalid
			VexRiscvAvalon_0_irq_controller_waitrequest        => mm_interconnect_0_vexriscvavalon_0_irq_controller_waitrequest    --                                             .waitrequest
		);

	mm_interconnect_1 : component qsys0_mm_interconnect_1
		port map (
			clk_0_clk_clk                                      => clk_clk,                                                        --                                    clk_0_clk.clk
			VexRiscvAvalon_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                 -- VexRiscvAvalon_0_reset_reset_bridge_in_reset.reset
			VexRiscvAvalon_0_instruction_bus_address           => vexriscvavalon_0_instruction_bus_address,                       --             VexRiscvAvalon_0_instruction_bus.address
			VexRiscvAvalon_0_instruction_bus_waitrequest       => mm_interconnect_1_vexriscvavalon_0_instruction_bus_waitrequest, --                                             .waitrequest
			VexRiscvAvalon_0_instruction_bus_read              => vexriscvavalon_0_instruction_bus_read,                          --                                             .read
			VexRiscvAvalon_0_instruction_bus_readdata          => vexriscvavalon_0_instruction_bus_readdata,                      --                                             .readdata
			VexRiscvAvalon_0_instruction_bus_readdatavalid     => vexriscvavalon_0_instruction_bus_readdatavalid,                 --                                             .readdatavalid
			VexRiscvAvalon_0_instruction_bus_response          => vexriscvavalon_0_instruction_bus_response,                      --                                             .response
			onchip_memory2_0_s1_address                        => mm_interconnect_1_onchip_memory2_0_s1_address,                  --                          onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                          => mm_interconnect_1_onchip_memory2_0_s1_write,                    --                                             .write
			onchip_memory2_0_s1_readdata                       => mm_interconnect_1_onchip_memory2_0_s1_readdata,                 --                                             .readdata
			onchip_memory2_0_s1_writedata                      => mm_interconnect_1_onchip_memory2_0_s1_writedata,                --                                             .writedata
			onchip_memory2_0_s1_byteenable                     => mm_interconnect_1_onchip_memory2_0_s1_byteenable,               --                                             .byteenable
			onchip_memory2_0_s1_chipselect                     => mm_interconnect_1_onchip_memory2_0_s1_chipselect,               --                                             .chipselect
			onchip_memory2_0_s1_clken                          => mm_interconnect_1_onchip_memory2_0_s1_clken                     --                                             .clken
		);

	irq_mapper : component qsys0_irq_mapper
		port map (
			clk           => clk_clk,                                 --       clk.clk
			reset         => rst_controller_reset_out_reset,          -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,                -- receiver0.irq
			sender_irq    => vexriscvavalon_0_interrupt_receiver_irq  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	vexriscvavalon_0_data_bus_inv <= not mm_interconnect_0_vexriscvavalon_0_data_bus_waitrequest;

	mm_interconnect_0_pio_0_s1_write_ports_inv <= not mm_interconnect_0_pio_0_s1_write;

	mm_interconnect_0_uart_0_s1_read_ports_inv <= not mm_interconnect_0_uart_0_s1_read;

	mm_interconnect_0_uart_0_s1_write_ports_inv <= not mm_interconnect_0_uart_0_s1_write;

	vexriscvavalon_0_instruction_bus_inv <= not mm_interconnect_1_vexriscvavalon_0_instruction_bus_waitrequest;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of qsys0
