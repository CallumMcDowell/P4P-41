-- vexriscv_system.vhd

-- Generated using ACDS version 21.1 850

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity vexriscv_system is
	port (
		clk_clk                                          : in  std_logic := '0'; --                                       clk.clk
		reset_reset_n                                    : in  std_logic := '0'; --                                     reset.reset_n
		vexriscvavalonmaxperf_0_jtag_tms                 : in  std_logic := '0'; --              vexriscvavalonmaxperf_0_jtag.tms
		vexriscvavalonmaxperf_0_jtag_tdi                 : in  std_logic := '0'; --                                          .tdi
		vexriscvavalonmaxperf_0_jtag_tdo                 : out std_logic;        --                                          .tdo
		vexriscvavalonmaxperf_0_jtag_tck                 : in  std_logic := '0'; --                                          .tck
		vexriscvavalonmaxperf_0_softwareinterrupt_export : in  std_logic := '0'  -- vexriscvavalonmaxperf_0_softwareinterrupt.export
	);
end entity vexriscv_system;

architecture rtl of vexriscv_system is
	component VexRiscvAvalonMaxPerf is
		port (
			timerInterrupt           : in  std_logic                     := 'X';             -- irq
			externalInterrupt        : in  std_logic                     := 'X';             -- irq
			softwareInterrupt        : in  std_logic                     := 'X';             -- export
			debug_resetOut           : out std_logic;                                        -- reset
			iBusAvalon_address       : out std_logic_vector(31 downto 0);                    -- address
			iBusAvalon_read          : out std_logic;                                        -- read
			iBusAvalon_waitRequestn  : in  std_logic                     := 'X';             -- waitrequest_n
			iBusAvalon_burstCount    : out std_logic_vector(3 downto 0);                     -- burstcount
			iBusAvalon_response      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			iBusAvalon_readDataValid : in  std_logic                     := 'X';             -- readdatavalid
			iBusAvalon_readData      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dBusAvalon_address       : out std_logic_vector(31 downto 0);                    -- address
			dBusAvalon_read          : out std_logic;                                        -- read
			dBusAvalon_write         : out std_logic;                                        -- write
			dBusAvalon_waitRequestn  : in  std_logic                     := 'X';             -- waitrequest_n
			dBusAvalon_burstCount    : out std_logic_vector(3 downto 0);                     -- burstcount
			dBusAvalon_byteEnable    : out std_logic_vector(3 downto 0);                     -- byteenable
			dBusAvalon_writeData     : out std_logic_vector(31 downto 0);                    -- writedata
			dBusAvalon_response      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			dBusAvalon_readDataValid : in  std_logic                     := 'X';             -- readdatavalid
			dBusAvalon_readData      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_tms                 : in  std_logic                     := 'X';             -- export
			jtag_tdi                 : in  std_logic                     := 'X';             -- export
			jtag_tdo                 : out std_logic;                                        -- export
			jtag_tck                 : in  std_logic                     := 'X';             -- export
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			debugReset               : in  std_logic                     := 'X'              -- reset
		);
	end component VexRiscvAvalonMaxPerf;

	component vexriscv_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component vexriscv_system_jtag_uart_0;

	component vexriscv_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                             : in  std_logic                     := 'X';             -- clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			VexRiscvAvalonMaxPerf_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			VexRiscvAvalonMaxPerf_0_dBusAvalon_address                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			VexRiscvAvalonMaxPerf_0_dBusAvalon_waitrequest            : out std_logic;                                        -- waitrequest
			VexRiscvAvalonMaxPerf_0_dBusAvalon_burstcount             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			VexRiscvAvalonMaxPerf_0_dBusAvalon_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			VexRiscvAvalonMaxPerf_0_dBusAvalon_read                   : in  std_logic                     := 'X';             -- read
			VexRiscvAvalonMaxPerf_0_dBusAvalon_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			VexRiscvAvalonMaxPerf_0_dBusAvalon_readdatavalid          : out std_logic;                                        -- readdatavalid
			VexRiscvAvalonMaxPerf_0_dBusAvalon_write                  : in  std_logic                     := 'X';             -- write
			VexRiscvAvalonMaxPerf_0_dBusAvalon_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			VexRiscvAvalonMaxPerf_0_dBusAvalon_response               : out std_logic_vector(1 downto 0);                     -- response
			VexRiscvAvalonMaxPerf_0_iBusAvalon_address                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			VexRiscvAvalonMaxPerf_0_iBusAvalon_waitrequest            : out std_logic;                                        -- waitrequest
			VexRiscvAvalonMaxPerf_0_iBusAvalon_burstcount             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			VexRiscvAvalonMaxPerf_0_iBusAvalon_read                   : in  std_logic                     := 'X';             -- read
			VexRiscvAvalonMaxPerf_0_iBusAvalon_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			VexRiscvAvalonMaxPerf_0_iBusAvalon_readdatavalid          : out std_logic;                                        -- readdatavalid
			VexRiscvAvalonMaxPerf_0_iBusAvalon_response               : out std_logic_vector(1 downto 0);                     -- response
			jtag_uart_0_avalon_jtag_slave_address                     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                       : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                        : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                  : out std_logic                                         -- chipselect
		);
	end component vexriscv_system_mm_interconnect_0;

	component vexriscv_system_irq_mapper is
		port (
			clk        : in  std_logic                    := 'X'; -- clk
			reset      : in  std_logic                    := 'X'; -- reset
			sender_irq : out std_logic_vector(0 downto 0)         -- irq
		);
	end component vexriscv_system_irq_mapper;

	component vexriscv_system_irq_mapper_001 is
		port (
			clk           : in  std_logic                    := 'X'; -- clk
			reset         : in  std_logic                    := 'X'; -- reset
			receiver0_irq : in  std_logic                    := 'X'; -- irq
			sender_irq    : out std_logic_vector(0 downto 0)         -- irq
		);
	end component vexriscv_system_irq_mapper_001;

	component vexriscv_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component vexriscv_system_rst_controller;

	component vexriscv_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component vexriscv_system_rst_controller_001;

	signal mm_interconnect_0_vexriscvavalonmaxperf_0_dbusavalon_waitrequest : std_logic;                     -- mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_waitrequest -> mm_interconnect_0_vexriscvavalonmaxperf_0_dbusavalon_waitrequest:in
	signal vexriscvavalonmaxperf_0_dbusavalon_readdata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_readdata -> VexRiscvAvalonMaxPerf_0:dBusAvalon_readData
	signal vexriscvavalonmaxperf_0_dbusavalon_address                       : std_logic_vector(31 downto 0); -- VexRiscvAvalonMaxPerf_0:dBusAvalon_address -> mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_address
	signal vexriscvavalonmaxperf_0_dbusavalon_read                          : std_logic;                     -- VexRiscvAvalonMaxPerf_0:dBusAvalon_read -> mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_read
	signal vexriscvavalonmaxperf_0_dbusavalon_byteenable                    : std_logic_vector(3 downto 0);  -- VexRiscvAvalonMaxPerf_0:dBusAvalon_byteEnable -> mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_byteenable
	signal vexriscvavalonmaxperf_0_dbusavalon_readdatavalid                 : std_logic;                     -- mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_readdatavalid -> VexRiscvAvalonMaxPerf_0:dBusAvalon_readDataValid
	signal vexriscvavalonmaxperf_0_dbusavalon_response                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_response -> VexRiscvAvalonMaxPerf_0:dBusAvalon_response
	signal vexriscvavalonmaxperf_0_dbusavalon_write                         : std_logic;                     -- VexRiscvAvalonMaxPerf_0:dBusAvalon_write -> mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_write
	signal vexriscvavalonmaxperf_0_dbusavalon_writedata                     : std_logic_vector(31 downto 0); -- VexRiscvAvalonMaxPerf_0:dBusAvalon_writeData -> mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_writedata
	signal vexriscvavalonmaxperf_0_dbusavalon_burstcount                    : std_logic_vector(3 downto 0);  -- VexRiscvAvalonMaxPerf_0:dBusAvalon_burstCount -> mm_interconnect_0:VexRiscvAvalonMaxPerf_0_dBusAvalon_burstcount
	signal mm_interconnect_0_vexriscvavalonmaxperf_0_ibusavalon_waitrequest : std_logic;                     -- mm_interconnect_0:VexRiscvAvalonMaxPerf_0_iBusAvalon_waitrequest -> mm_interconnect_0_vexriscvavalonmaxperf_0_ibusavalon_waitrequest:in
	signal vexriscvavalonmaxperf_0_ibusavalon_readdata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:VexRiscvAvalonMaxPerf_0_iBusAvalon_readdata -> VexRiscvAvalonMaxPerf_0:iBusAvalon_readData
	signal vexriscvavalonmaxperf_0_ibusavalon_address                       : std_logic_vector(31 downto 0); -- VexRiscvAvalonMaxPerf_0:iBusAvalon_address -> mm_interconnect_0:VexRiscvAvalonMaxPerf_0_iBusAvalon_address
	signal vexriscvavalonmaxperf_0_ibusavalon_read                          : std_logic;                     -- VexRiscvAvalonMaxPerf_0:iBusAvalon_read -> mm_interconnect_0:VexRiscvAvalonMaxPerf_0_iBusAvalon_read
	signal vexriscvavalonmaxperf_0_ibusavalon_readdatavalid                 : std_logic;                     -- mm_interconnect_0:VexRiscvAvalonMaxPerf_0_iBusAvalon_readdatavalid -> VexRiscvAvalonMaxPerf_0:iBusAvalon_readDataValid
	signal vexriscvavalonmaxperf_0_ibusavalon_response                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:VexRiscvAvalonMaxPerf_0_iBusAvalon_response -> VexRiscvAvalonMaxPerf_0:iBusAvalon_response
	signal vexriscvavalonmaxperf_0_ibusavalon_burstcount                    : std_logic_vector(3 downto 0);  -- VexRiscvAvalonMaxPerf_0:iBusAvalon_burstCount -> mm_interconnect_0:VexRiscvAvalonMaxPerf_0_iBusAvalon_burstcount
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect       : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata         : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest      : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read             : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal vexriscvavalonmaxperf_0_timerinterrupt_irq                       : std_logic;                     -- irq_mapper:sender_irq -> VexRiscvAvalonMaxPerf_0:timerInterrupt
	signal irq_mapper_001_receiver0_irq                                     : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper_001:receiver0_irq
	signal vexriscvavalonmaxperf_0_externalinterrupt_irq                    : std_logic;                     -- irq_mapper_001:sender_irq -> VexRiscvAvalonMaxPerf_0:externalInterrupt
	signal rst_controller_reset_out_reset                                   : std_logic;                     -- rst_controller:reset_out -> [VexRiscvAvalonMaxPerf_0:reset, irq_mapper:reset, irq_mapper_001:reset, mm_interconnect_0:VexRiscvAvalonMaxPerf_0_reset_reset_bridge_in_reset_reset]
	signal vexriscvavalonmaxperf_0_debug_resetout_reset                     : std_logic;                     -- VexRiscvAvalonMaxPerf_0:debug_resetOut -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset                               : std_logic;                     -- rst_controller_001:reset_out -> [VexRiscvAvalonMaxPerf_0:debugReset, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                          : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal vexriscvavalonmaxperf_0_dbusavalon_inv                           : std_logic;                     -- mm_interconnect_0_vexriscvavalonmaxperf_0_dbusavalon_waitrequest:inv -> VexRiscvAvalonMaxPerf_0:dBusAvalon_waitRequestn
	signal vexriscvavalonmaxperf_0_ibusavalon_inv                           : std_logic;                     -- mm_interconnect_0_vexriscvavalonmaxperf_0_ibusavalon_waitrequest:inv -> VexRiscvAvalonMaxPerf_0:iBusAvalon_waitRequestn
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv   : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal rst_controller_001_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> jtag_uart_0:rst_n

begin

	vexriscvavalonmaxperf_0 : component VexRiscvAvalonMaxPerf
		port map (
			timerInterrupt           => vexriscvavalonmaxperf_0_timerinterrupt_irq,       --    timerInterrupt.irq
			externalInterrupt        => vexriscvavalonmaxperf_0_externalinterrupt_irq,    -- externalInterrupt.irq
			softwareInterrupt        => vexriscvavalonmaxperf_0_softwareinterrupt_export, -- softwareInterrupt.export
			debug_resetOut           => vexriscvavalonmaxperf_0_debug_resetout_reset,     --    debug_resetOut.reset
			iBusAvalon_address       => vexriscvavalonmaxperf_0_ibusavalon_address,       --        iBusAvalon.address
			iBusAvalon_read          => vexriscvavalonmaxperf_0_ibusavalon_read,          --                  .read
			iBusAvalon_waitRequestn  => vexriscvavalonmaxperf_0_ibusavalon_inv,           --                  .waitrequest_n
			iBusAvalon_burstCount    => vexriscvavalonmaxperf_0_ibusavalon_burstcount,    --                  .burstcount
			iBusAvalon_response      => vexriscvavalonmaxperf_0_ibusavalon_response,      --                  .response
			iBusAvalon_readDataValid => vexriscvavalonmaxperf_0_ibusavalon_readdatavalid, --                  .readdatavalid
			iBusAvalon_readData      => vexriscvavalonmaxperf_0_ibusavalon_readdata,      --                  .readdata
			dBusAvalon_address       => vexriscvavalonmaxperf_0_dbusavalon_address,       --        dBusAvalon.address
			dBusAvalon_read          => vexriscvavalonmaxperf_0_dbusavalon_read,          --                  .read
			dBusAvalon_write         => vexriscvavalonmaxperf_0_dbusavalon_write,         --                  .write
			dBusAvalon_waitRequestn  => vexriscvavalonmaxperf_0_dbusavalon_inv,           --                  .waitrequest_n
			dBusAvalon_burstCount    => vexriscvavalonmaxperf_0_dbusavalon_burstcount,    --                  .burstcount
			dBusAvalon_byteEnable    => vexriscvavalonmaxperf_0_dbusavalon_byteenable,    --                  .byteenable
			dBusAvalon_writeData     => vexriscvavalonmaxperf_0_dbusavalon_writedata,     --                  .writedata
			dBusAvalon_response      => vexriscvavalonmaxperf_0_dbusavalon_response,      --                  .response
			dBusAvalon_readDataValid => vexriscvavalonmaxperf_0_dbusavalon_readdatavalid, --                  .readdatavalid
			dBusAvalon_readData      => vexriscvavalonmaxperf_0_dbusavalon_readdata,      --                  .readdata
			jtag_tms                 => vexriscvavalonmaxperf_0_jtag_tms,                 --              jtag.export
			jtag_tdi                 => vexriscvavalonmaxperf_0_jtag_tdi,                 --                  .export
			jtag_tdo                 => vexriscvavalonmaxperf_0_jtag_tdo,                 --                  .export
			jtag_tck                 => vexriscvavalonmaxperf_0_jtag_tck,                 --                  .export
			clk                      => clk_clk,                                          --               clk.clk
			reset                    => rst_controller_reset_out_reset,                   --             reset.reset
			debugReset               => rst_controller_001_reset_out_reset                --        debugReset.reset
		);

	jtag_uart_0 : component vexriscv_system_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver0_irq                                     --               irq.irq
		);

	mm_interconnect_0 : component vexriscv_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                             => clk_clk,                                                          --                                           clk_0_clk.clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset             => rst_controller_001_reset_out_reset,                               --             jtag_uart_0_reset_reset_bridge_in_reset.reset
			VexRiscvAvalonMaxPerf_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                   -- VexRiscvAvalonMaxPerf_0_reset_reset_bridge_in_reset.reset
			VexRiscvAvalonMaxPerf_0_dBusAvalon_address                => vexriscvavalonmaxperf_0_dbusavalon_address,                       --                  VexRiscvAvalonMaxPerf_0_dBusAvalon.address
			VexRiscvAvalonMaxPerf_0_dBusAvalon_waitrequest            => mm_interconnect_0_vexriscvavalonmaxperf_0_dbusavalon_waitrequest, --                                                    .waitrequest
			VexRiscvAvalonMaxPerf_0_dBusAvalon_burstcount             => vexriscvavalonmaxperf_0_dbusavalon_burstcount,                    --                                                    .burstcount
			VexRiscvAvalonMaxPerf_0_dBusAvalon_byteenable             => vexriscvavalonmaxperf_0_dbusavalon_byteenable,                    --                                                    .byteenable
			VexRiscvAvalonMaxPerf_0_dBusAvalon_read                   => vexriscvavalonmaxperf_0_dbusavalon_read,                          --                                                    .read
			VexRiscvAvalonMaxPerf_0_dBusAvalon_readdata               => vexriscvavalonmaxperf_0_dbusavalon_readdata,                      --                                                    .readdata
			VexRiscvAvalonMaxPerf_0_dBusAvalon_readdatavalid          => vexriscvavalonmaxperf_0_dbusavalon_readdatavalid,                 --                                                    .readdatavalid
			VexRiscvAvalonMaxPerf_0_dBusAvalon_write                  => vexriscvavalonmaxperf_0_dbusavalon_write,                         --                                                    .write
			VexRiscvAvalonMaxPerf_0_dBusAvalon_writedata              => vexriscvavalonmaxperf_0_dbusavalon_writedata,                     --                                                    .writedata
			VexRiscvAvalonMaxPerf_0_dBusAvalon_response               => vexriscvavalonmaxperf_0_dbusavalon_response,                      --                                                    .response
			VexRiscvAvalonMaxPerf_0_iBusAvalon_address                => vexriscvavalonmaxperf_0_ibusavalon_address,                       --                  VexRiscvAvalonMaxPerf_0_iBusAvalon.address
			VexRiscvAvalonMaxPerf_0_iBusAvalon_waitrequest            => mm_interconnect_0_vexriscvavalonmaxperf_0_ibusavalon_waitrequest, --                                                    .waitrequest
			VexRiscvAvalonMaxPerf_0_iBusAvalon_burstcount             => vexriscvavalonmaxperf_0_ibusavalon_burstcount,                    --                                                    .burstcount
			VexRiscvAvalonMaxPerf_0_iBusAvalon_read                   => vexriscvavalonmaxperf_0_ibusavalon_read,                          --                                                    .read
			VexRiscvAvalonMaxPerf_0_iBusAvalon_readdata               => vexriscvavalonmaxperf_0_ibusavalon_readdata,                      --                                                    .readdata
			VexRiscvAvalonMaxPerf_0_iBusAvalon_readdatavalid          => vexriscvavalonmaxperf_0_ibusavalon_readdatavalid,                 --                                                    .readdatavalid
			VexRiscvAvalonMaxPerf_0_iBusAvalon_response               => vexriscvavalonmaxperf_0_ibusavalon_response,                      --                                                    .response
			jtag_uart_0_avalon_jtag_slave_address                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,          --                       jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,            --                                                    .write
			jtag_uart_0_avalon_jtag_slave_read                        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,             --                                                    .read
			jtag_uart_0_avalon_jtag_slave_readdata                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,         --                                                    .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,        --                                                    .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,      --                                                    .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect        --                                                    .chipselect
		);

	irq_mapper : component vexriscv_system_irq_mapper
		port map (
			clk           => clk_clk,                                    --       clk.clk
			reset         => rst_controller_reset_out_reset,             -- clk_reset.reset
			sender_irq(0) => vexriscvavalonmaxperf_0_timerinterrupt_irq  --    sender.irq
		);

	irq_mapper_001 : component vexriscv_system_irq_mapper_001
		port map (
			clk           => clk_clk,                                       --       clk.clk
			reset         => rst_controller_reset_out_reset,                -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq,                  -- receiver0.irq
			sender_irq(0) => vexriscvavalonmaxperf_0_externalinterrupt_irq  --    sender.irq
		);

	rst_controller : component vexriscv_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                      -- reset_in0.reset
			reset_in1      => vexriscvavalonmaxperf_0_debug_resetout_reset, -- reset_in1.reset
			clk            => clk_clk,                                      --       clk.clk
			reset_out      => rst_controller_reset_out_reset,               -- reset_out.reset
			reset_req      => open,                                         -- (terminated)
			reset_req_in0  => '0',                                          -- (terminated)
			reset_req_in1  => '0',                                          -- (terminated)
			reset_in2      => '0',                                          -- (terminated)
			reset_req_in2  => '0',                                          -- (terminated)
			reset_in3      => '0',                                          -- (terminated)
			reset_req_in3  => '0',                                          -- (terminated)
			reset_in4      => '0',                                          -- (terminated)
			reset_req_in4  => '0',                                          -- (terminated)
			reset_in5      => '0',                                          -- (terminated)
			reset_req_in5  => '0',                                          -- (terminated)
			reset_in6      => '0',                                          -- (terminated)
			reset_req_in6  => '0',                                          -- (terminated)
			reset_in7      => '0',                                          -- (terminated)
			reset_req_in7  => '0',                                          -- (terminated)
			reset_in8      => '0',                                          -- (terminated)
			reset_req_in8  => '0',                                          -- (terminated)
			reset_in9      => '0',                                          -- (terminated)
			reset_req_in9  => '0',                                          -- (terminated)
			reset_in10     => '0',                                          -- (terminated)
			reset_req_in10 => '0',                                          -- (terminated)
			reset_in11     => '0',                                          -- (terminated)
			reset_req_in11 => '0',                                          -- (terminated)
			reset_in12     => '0',                                          -- (terminated)
			reset_req_in12 => '0',                                          -- (terminated)
			reset_in13     => '0',                                          -- (terminated)
			reset_req_in13 => '0',                                          -- (terminated)
			reset_in14     => '0',                                          -- (terminated)
			reset_req_in14 => '0',                                          -- (terminated)
			reset_in15     => '0',                                          -- (terminated)
			reset_req_in15 => '0'                                           -- (terminated)
		);

	rst_controller_001 : component vexriscv_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	vexriscvavalonmaxperf_0_dbusavalon_inv <= not mm_interconnect_0_vexriscvavalonmaxperf_0_dbusavalon_waitrequest;

	vexriscvavalonmaxperf_0_ibusavalon_inv <= not mm_interconnect_0_vexriscvavalonmaxperf_0_ibusavalon_waitrequest;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of vexriscv_system
